module main

import cjson  // import lydiandy.cjson


fn main() {
	// print json 
	user := cjson.obj()
	user.set("name", cjson.str("Tom"))
	user.set("age", cjson.num(18))
	user.set("gender", cjson.boolean(true))
	user.set("password", cjson.null())

	friends := cjson.list()
	friend := cjson.obj()
	friend.set("name", cjson.str("Jack"))
	friends.add(friend)
	user.set("friends", friends)

	leader := cjson.obj()
	leader.set("name", cjson.str("Mike"))
	user.set('leader', leader)

	json_str := user.dump()
	println(json_str)

	// parse json 
	json_content:='{"name":"jack","age":22}'
	res:=cjson.json_parse(json_content)

	// {
    //     "name": "Tom",
    //     "age":  18,
    //     "gender":       true,
    //     "password":     null,
    //     "friends":      [{
    //                     "name": "Jack"
    //             }],
    //     "leader":       {
    //             "name": "Mike"
    //     }
	// }
	
	name:=cjson.get_object_item(res,'name')
	age:=cjson.get_object_item(res,'age')
	println(name.valuestring)
	println(age.valueint)
}
